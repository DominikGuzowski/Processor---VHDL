----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 26.12.2020 18:00:12
-- Design Name: 
-- Module Name: Memory2p9_32Bit - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Memory2p9_32Bit is
    Port ( Address : in STD_LOGIC_VECTOR (31 downto 0);
           MW : in STD_LOGIC;
           Clk : in STD_LOGIC;
           Data_in : in STD_LOGIC_VECTOR (31 downto 0);
           Data_out : out STD_LOGIC_VECTOR (31 downto 0));
end Memory2p9_32Bit;
--MW 0 allows to read data, MW 1 allows to write data.
architecture Behavioral of Memory2p9_32Bit is
type Mem_Array is array(0 to 511) of std_logic_vector(31 downto 0);
constant DELAY : Time := 5ns;
constant INIT_0 : std_logic_vector(7 downto 0) := x"07"; --Loads 0 into registers 0-31 (SHOULD NOT BE USED BY PROGRAMMER)
constant INIT_1 : std_logic_vector(7 downto 0) := x"01"; --Loads 0 into register 32 (SHOULD NOT BE USER BY PROGRAMMER)
constant IN_SKP : std_logic_vector(7 downto 0) := x"08"; --Skips 1 clock cycle.
constant IN_AND : std_logic_vector(7 downto 0) := x"0A"; --INSTRUCTION: And 
constant IN_ORR : std_logic_vector(7 downto 0) := x"0B"; --INSTRUCTION: Or
constant IN_XOR : std_logic_vector(7 downto 0) := x"0C"; --INSTRUCTION: Xor
constant IN_NOT : std_logic_vector(7 downto 0) := x"0D"; --INSTRUCTION: Not
constant IN_MVI : std_logic_vector(7 downto 0) := x"0E"; --INSTRUCTION: Move immediate (5 bit)
constant IN_MOV : std_logic_vector(7 downto 0) := x"0F"; --INSTRUCTION: Move
constant IN_ADD : std_logic_vector(7 downto 0) := x"10"; --INSTRUCTION: Add
constant IN_ADI : std_logic_vector(7 downto 0) := x"11"; --INSTRUCTION: Add immediate (5 bit)
constant IN_INC : std_logic_vector(7 downto 0) := x"12"; --INSTRUCTION: Increment
constant IN_ADC : std_logic_vector(7 downto 0) := x"13"; --INSTRUCTION: Add with Carry
constant IN_AOC : std_logic_vector(7 downto 0) := x"14"; --INSTRUCTION: Add with 1s Compliment of R[SB]
constant IN_SUB : std_logic_vector(7 downto 0) := x"15"; --INSTRUCTION: Subtract
constant IN_SBI : std_logic_vector(7 downto 0) := x"16"; --INSTRUCTION: Subtract immediate (5 bit)
constant IN_DEC : std_logic_vector(7 downto 0) := x"17"; --INSTRUCTION: Decrement
constant IN_LDR : std_logic_vector(7 downto 0) := x"18"; --INSTRUCTION: Load Register
constant IN_LSL : std_logic_vector(7 downto 0) := x"1A"; --INSTRUCTION: Logical Shift Left
constant IN_LSR : std_logic_vector(7 downto 0) := x"1B"; --INSTRUCTION: Logical Shift Right
constant IN_STR : std_logic_vector(7 downto 0) := x"1C"; --INSTRUCTION: Store Register
constant IN_SRM : std_logic_vector(7 downto 0) := x"20"; --INSTRUCTION: Logical shift right multiple times (defined by #N)
constant IN_SLM : std_logic_vector(7 downto 0) := x"28"; --INSTRUCTION: Logical shift left multiple times (defined by #N)
constant IN_BAL : std_logic_vector(7 downto 0) := x"30"; --INSTRUCTION: Branch always
constant IN_BNS : std_logic_vector(7 downto 0) := x"33"; --INSTRUCTION: Branch if N set
constant IN_BZS : std_logic_vector(7 downto 0) := x"35"; --INSTRUCTION: Branch if Z set
constant IN_BVS : std_logic_vector(7 downto 0) := x"37"; --INSTRUCTION: Branch if V set
constant IN_BCS : std_logic_vector(7 downto 0) := x"39"; --INSTRUCTION: Branch if C set
constant IN_BZC : std_logic_vector(7 downto 0) := x"3B"; --INSTRUCTION: Branch if Z clear
constant IN_BCC : std_logic_vector(7 downto 0) := x"3D"; --INSTRUCTION: Branch if C clear
constant IN_CMP : std_logic_vector(7 downto 0) := x"40"; --INSTRUCTION: Compare
constant IN_CPI : std_logic_vector(7 downto 0) := x"41"; --INSTRUCTION: Compare immediate (5 bits)
constant IN_BEQ : std_logic_vector(7 downto 0) := x"42"; --INSTRUCTION: Branch if a == b
constant IN_BNE : std_logic_vector(7 downto 0) := x"44"; --INSTRUCTION: Branch if a != b
constant IN_BHS : std_logic_vector(7 downto 0) := x"46"; --INSTRUCTION: Branch if a >= b (unsigned)
constant IN_BLO : std_logic_vector(7 downto 0) := x"48"; --INSTRUCTION: Branch if a < b (unsigned)
constant IN_BPL : std_logic_vector(7 downto 0) := x"4A"; --INSTRUCTION: Branch if a >= 0
constant IN_BMI : std_logic_vector(7 downto 0) := x"4C"; --INSTRUCTION: Branch if a < 0
constant IN_BHI : std_logic_vector(7 downto 0) := x"4E"; --INSTRUCTION: Branch if a > b (unsigned)
constant IN_BLS : std_logic_vector(7 downto 0) := x"51"; --INSTRUCTION: Branch if a <= b (unsigned)
constant IN_BGE : std_logic_vector(7 downto 0) := x"54"; --INSTRUCTION: Branch if a >= b
constant IN_BLT : std_logic_vector(7 downto 0) := x"59"; --INSTRUCTION: Branch if a < b
constant IN_BGT : std_logic_vector(7 downto 0) := x"5E"; --INSTRUCTION: Branch if a > b
constant IN_BLE : std_logic_vector(7 downto 0) := x"60"; --INSTRUCTION: Branch if a <= b
constant IN_END : std_logic_vector(7 downto 0) := x"02"; --INSTRUCTION: Ends the program.
constant NO_INS : std_logic_vector(7 downto 0) := x"05"; --No instruction        
begin
Mem_Process: process(Address, Data_in, Clk)
variable Mem_Data : Mem_Array := (
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & INIT_0 & "00000" & "00000" & "00000", --0x00
 "000000000" & INIT_0 & "00001" & "00000" & "00000", --0x01
 "000000000" & INIT_0 & "00010" & "00000" & "00000", --0x02
 "000000000" & INIT_0 & "00011" & "00000" & "00000", --0x03
 "000000000" & INIT_0 & "00100" & "00000" & "00000", --0x04
 "000000000" & INIT_0 & "00101" & "00000" & "00000", --0x05
 "000000000" & INIT_0 & "00110" & "00000" & "00000", --0x06
 "000000000" & INIT_0 & "00111" & "00000" & "00000", --0x07
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & INIT_0 & "01000" & "00000" & "00000", --0x08
 "000000000" & INIT_0 & "01001" & "00000" & "00000", --0x09
 "000000000" & INIT_0 & "01010" & "00000" & "00000", --0x0A
 "000000000" & INIT_0 & "01011" & "00000" & "00000", --0x0B
 "000000000" & INIT_0 & "01100" & "00000" & "00000", --0x0C
 "000000000" & INIT_0 & "01101" & "00000" & "00000", --0x0D
 "000000000" & INIT_0 & "01110" & "00000" & "00000", --0x0E
 "000000000" & INIT_0 & "01111" & "00000" & "00000", --0x0F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & INIT_0 & "10000" & "00000" & "00000", --0x10
 "000000000" & INIT_0 & "10001" & "00000" & "00000", --0x11
 "000000000" & INIT_0 & "10010" & "00000" & "00000", --0x12
 "000000000" & INIT_0 & "10011" & "00000" & "00000", --0x13
 "000000000" & INIT_0 & "10100" & "00000" & "00000", --0x14
 "000000000" & INIT_0 & "10101" & "00000" & "00000", --0x15
 "000000000" & INIT_0 & "10110" & "00000" & "00000", --0x16
 "000000000" & INIT_0 & "10111" & "00000" & "00000", --0x17
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & INIT_0 & "11000" & "00000" & "00000", --0x18
 "000000000" & INIT_0 & "11001" & "00000" & "00000", --0x19
 "000000000" & INIT_0 & "11010" & "00000" & "00000", --0x1A
 "000000000" & INIT_0 & "11011" & "00000" & "00000", --0x1B
 "000000000" & INIT_0 & "11100" & "00000" & "00000", --0x1C
 "000000000" & INIT_0 & "11101" & "00000" & "00000", --0x1D
 "000000000" & INIT_0 & "11110" & "00000" & "00000", --0x1E
 "000000000" & INIT_1 & "11111" & "00000" & "00000", --0x1F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |          END OF INITIALIZATION: First instruction fetch goes on line 0x20
 "000000000" & IN_MVI & "00000" & "00000" & "00000", --0x20 FETCH MVI
 "000000000" & IN_ADD & "00000" & "00000" & "10000", --0x21 FETCH ADD DECODE MVI
 "000000000" & IN_ADD & "00000" & "00000" & "00000", --0x22 FETCH ADD DECODE ADD EXECUTE MVI
 "000000000" & IN_LDR & "00000" & "00000" & "00000", --0x23 FETCH LDR DECODE ADD EXECUTE ADD
 "000000000" & IN_MVI & "00001" & "00000" & "00000", --0x24 FETCH MVI DECODE LDR EXECUTE ADD
 "000000000" & IN_STR & "00010" & "00000" & "00001", --0x25 FETCH STR DECODE MVI EXECUTE LDR
 "000000000" & IN_LDR & "00000" & "00000" & "00010", --0x26 FETCH LDR DECODE STR EXECUTE MVI
 "000000000" & IN_CMP & "00011" & "00000" & "00000", --0x27 FETCH CMP DECODE LDR EXECUTE STR
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB 
 "000000000" & IN_BGT & "00000" & "00010" & "00001", --0x28 FETCH BGT DECODE CMP EXECUTE LDR
 "000000000" & IN_MVI & "00000" & "00000" & "00011", --0x29 FETCH MVI DECODE BGT EXECUTE CMP <-Set OFFSET
 "000000000" & IN_END & "00101" & "00000" & "01111", --0x2A FETCH END DECODE MVI EXECUTE BGT
 "000000000" & NO_INS & "00000" & "00000" & "00000", --0x2B FETCH --- DECODE END EXECUTE MVI
 "000000000" & NO_INS & "00000" & "00000" & "00000", --0x2C FETCH --- DECODE --- EXECUTE END
 "000000000" & IN_MVI & "00000" & "00000" & "00000", --0x2D FETCH MVI DECODE --- EXECUTE ---
 "000000000" & IN_INC & "00101" & "00000" & "01010", --0x2E FETCH END DECODE MVI EXECUTE ---
 "000000000" & IN_DEC & "00100" & "00100" & "00000", --0x2F  FETCH --- DECODE END EXECUTE MVI
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB   |
 "000000000" & IN_CPI & "00101" & "00101" & "00000", --0x30  FETCH --- DECODE --- EXECUTE END
 "000000000" & IN_BNE & "00000" & "00101" & "00000", --0x31  
 "000000000" & IN_ADI & "11111" & "00000" & "11011", --0x32 
 "000000000" & x"68" & "00100" & "00100" & "00110", --0x33 
 "000000000" & IN_END & "00100" & "00100" & "00101", --0x34 
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x35 
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x36 
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x37 
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x38 
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x39 
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x3A 
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x3B 
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x3C 
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x3D 
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x3E 
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x3F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "111111111" & x"FF" & "11111" & "11111" & "11111", --0x40 VALUE: -1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x41
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x42
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x43
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x44
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x45
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x46
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x47
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x48
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x49
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x4A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x4B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x4C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x4D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x4E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x4F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x50
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x51
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x52
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x53
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x54
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x55
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x56
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x57
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x58
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x59
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x5A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x5B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x5C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x5D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x5E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x5F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x60
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x61
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x62
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x63
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x64
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x65
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x66
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x67
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x68
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x69
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x6A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x6B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x6C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x6D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x6E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x6F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x70
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x71
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x72
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x73
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x74
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x75
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x76
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x77
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x78
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x79
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x7A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x7B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x7C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x7D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x7E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x7F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x80
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x81
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x82
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x83
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x84
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x85
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x86
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x87
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x88
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x89
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x8A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x8B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x8C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x8D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x8E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x8F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x90
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x91
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x92
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x93
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x94
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x95
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x96
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x97
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x98
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x99
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x9A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x9B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x9C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x9D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x9E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x9F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xA0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xA1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xA2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xA3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xA4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xA5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xA6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xA7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xA8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xA9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xAA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xAB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xAC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xAD
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xAE
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xAF
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xB0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xB1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xB2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xB3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xB4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xB5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xB6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xB7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xB8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xB9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xBA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xBB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xBC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xBD
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xBE
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xBF
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xC0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xC1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xC2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xC3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xC4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xC5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xC6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xC7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xC8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xC9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xCA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xCB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xCC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xCD
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xCE
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xCF
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xD0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xD1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xD2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xD3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xD4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xD5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xD6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xD7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xD8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xD9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xDA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xDB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xDC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xDD
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xDE
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xDF
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xE0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xE1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xE2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xE3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xE4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xE5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xE6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xE7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xE8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xE9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xEA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xEB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xEC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xED
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xEE
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xEF
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xF0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xF1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xF2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xF3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xF4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xF5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xF6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xF7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xF8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xF9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xFA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xFB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xFC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xFD
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xFE
 "000000000" & x"00" & "00000" & "00000" & "00000", --0xFF
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x100
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x101
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x102
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x103
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x104
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x105
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x106
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x107
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x108
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x109
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x10A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x10B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x10C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x10D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x10E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x10F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x110
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x111
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x112
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x113
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x114
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x115
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x116
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x117
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x118
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x119
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x11A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x11B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x11C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x11D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x11E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x11F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x120
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x121
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x122
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x123
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x124
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x125
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x126
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x127
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x128
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x129
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x12A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x12B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x12C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x12D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x12E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x12F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x130
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x131
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x132
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x133
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x134
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x135
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x136
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x137
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x138
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x139
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x13A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x13B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x13C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x13D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x13E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x13F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x140
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x141
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x142
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x143
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x144
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x145
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x146
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x147
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x148
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x149
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x14A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x14B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x14C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x14D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x14E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x14F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x150
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x151
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x152
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x153
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x154
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x155
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x156
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x157
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x158
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x159
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x15A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x15B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x15C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x15D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x15E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x15F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x160
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x161
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x162
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x163
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x164
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x165
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x166
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x167
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x168
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x169
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x16A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x16B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x16C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x16D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x16E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x16F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x170
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x171
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x172
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x173
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x174
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x175
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x176
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x177
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x178
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x179
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x17A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x17B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x17C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x17D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x17E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x17F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x180
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x181
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x182
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x183
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x184
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x185
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x186
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x187
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x188
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x189
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x18A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x18B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x18C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x18D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x18E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x18F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x190
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x191
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x192
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x193
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x194
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x195
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x196
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x197
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x198
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x199
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x19A
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x19B
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x19C
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x19D
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x19E
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x19F
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1A0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1A1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1A2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1A3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1A4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1A5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1A6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1A7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1A8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1A9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1AA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1AB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1AC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1AD
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1AE
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1AF
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1B0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1B1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1B2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1B3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1B4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1B5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1B6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1B7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1B8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1B9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1BA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1BB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1BC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1BD
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1BE
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1BF
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1C0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1C1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1C2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1C3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1C4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1C5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1C6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1C7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1C8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1C9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1CA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1CB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1CC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1CD
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1CE
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1CF
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1D0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1D1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1D2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1D3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1D4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1D5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1D6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1D7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1D8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1D9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1DA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1DB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1DC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1DD
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1DE
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1DF
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1E0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1E1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1E2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1E3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1E4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1E5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1E6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1E7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1E8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1E9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1EA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1EB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1EC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1ED
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1EE
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1EF
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1F0
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1F1
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1F2
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1F3
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1F4
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1F5
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1F6
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1F7
--|NOT USED| |Opcode|  | DR  |   | SA  |   | SB  |
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1F8
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1F9
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1FA
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1FB
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1FC
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1FD
 "000000000" & x"00" & "00000" & "00000" & "00000", --0x1FE
 "000000000" & x"00" & "00000" & "00000" & "00000"  --0x1FF
);
variable Adr : integer;
begin
Adr := conv_integer(unsigned(Address(8 downto 0)));
if MW = '1' and rising_edge(Clk) then
    Mem_Data(Adr) := Data_in;
end if;
Data_out <= Mem_Data(Adr) after DELAY;
end process;
end Behavioral;
